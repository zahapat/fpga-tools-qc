    -- Constants that are visible to all source files

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    package const_pack is

        constant QUBITS_CNT : natural := 4;
        -- constant QUBITS_CNT : natural := 6;
        -- constant QUBITS_CNT : natural := 8;
        
    end package;

    package body const_pack is

    end package body;