-- generics.vhd: This is an automatically generated file with generic parameters 
-- after running 'make generics' command.
package generics is

    constant INT_EMULATE_INPUTS : integer := 0;
    constant INT_QUBITS_CNT : integer := 4;
    constant INT_WHOLE_PHOTON_2H_DELAY_NS : integer := -2117;
    constant INT_DECIM_PHOTON_2H_DELAY_NS : integer := 95;
    constant INT_WHOLE_PHOTON_2V_DELAY_NS : integer := -2125;
    constant INT_DECIM_PHOTON_2V_DELAY_NS : integer := 35;
    constant INT_WHOLE_PHOTON_3H_DELAY_NS : integer := -1030;
    constant INT_DECIM_PHOTON_3H_DELAY_NS : integer := 35;
    constant INT_WHOLE_PHOTON_3V_DELAY_NS : integer := -1034;
    constant INT_DECIM_PHOTON_3V_DELAY_NS : integer := 45;
    constant INT_WHOLE_PHOTON_4H_DELAY_NS : integer := -3177;
    constant INT_DECIM_PHOTON_4H_DELAY_NS : integer := 95;
    constant INT_WHOLE_PHOTON_4V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_4V_DELAY_NS : integer := 05;
    constant INT_WHOLE_PHOTON_5H_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_5H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_5V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_5V_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_6H_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_6H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_6V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_6V_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_7H_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_7H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_7V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_7V_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_8H_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_8H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_8V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_8V_DELAY_NS : integer := 1;

end package generics;



package body generics is 

end package body generics;