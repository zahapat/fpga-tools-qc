    -- Signals that are visible to all source files

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    library lib_src;
    use lib_src.const_pack.all;
    use lib_src.types_pack.all;
    use lib_src.generics.all;

    package signals_pack is
        
    end package;

    package body signals_pack is

    end package body;