-- essentials_tb.vhd: This is an automatically generated file with information about 
-- project name and root directory after running 'make generics' command.
package essentials_tb is

    constant PROJ_NAME : string := "fpga-tools-qc";
    constant PROJ_DIR : string := "C:/Git/zahapat/fpga-tools-qc/";
    constant RANDOM_SEED_1 : natural := 1684619324;
    constant RANDOM_SEED_2 : natural := 787585433;

end package essentials_tb;



package body essentials_tb is 

end package body essentials_tb;