-- generics.vhd: This is an automatically generated file with generic parameters 
-- after running 'make generics' command.
package generics is

    constant INT_EMULATE_INPUTS : integer := 1;
    constant INT_QUBITS_CNT : integer := 4;
    constant INT_WHOLE_PHOTON_1H_DELAY_NS : integer := 75;
    constant INT_DECIM_PHOTON_1H_DELAY_NS : integer := 65;
    constant INT_WHOLE_PHOTON_1V_DELAY_NS : integer := 75;
    constant INT_DECIM_PHOTON_1V_DELAY_NS : integer := 01;
    constant INT_WHOLE_PHOTON_2H_DELAY_NS : integer := -1030;
    constant INT_DECIM_PHOTON_2H_DELAY_NS : integer := 95;
    constant INT_WHOLE_PHOTON_2V_DELAY_NS : integer := -1034;
    constant INT_DECIM_PHOTON_2V_DELAY_NS : integer := 35;
    constant INT_WHOLE_PHOTON_3H_DELAY_NS : integer := -2117;
    constant INT_DECIM_PHOTON_3H_DELAY_NS : integer := 35;
    constant INT_WHOLE_PHOTON_3V_DELAY_NS : integer := -2125;
    constant INT_DECIM_PHOTON_3V_DELAY_NS : integer := 45;
    constant INT_WHOLE_PHOTON_4H_DELAY_NS : integer := -3177;
    constant INT_DECIM_PHOTON_4H_DELAY_NS : integer := 95;
    constant INT_WHOLE_PHOTON_4V_DELAY_NS : integer := -3181;
    constant INT_DECIM_PHOTON_4V_DELAY_NS : integer := 0;
    constant INT_WHOLE_PHOTON_5H_DELAY_NS : integer := -4177;
    constant INT_DECIM_PHOTON_5H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_5V_DELAY_NS : integer := -4181;
    constant INT_DECIM_PHOTON_5V_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_6H_DELAY_NS : integer := -5177;
    constant INT_DECIM_PHOTON_6H_DELAY_NS : integer := 1;
    constant INT_WHOLE_PHOTON_6V_DELAY_NS : integer := -5181;
    constant INT_DECIM_PHOTON_6V_DELAY_NS : integer := 1;
    constant INT_CTRL_PULSE_HIGH_DURATION_NS : integer := 100;
    constant INT_CTRL_PULSE_DEAD_DURATION_NS : integer := 50;
    constant INT_CTRL_PULSE_EXTRA_DELAY_NS : integer := 0;
    constant INT_DISCARD_QUBITS_TIME_NS : integer := 0;

end package generics;



package body generics is 

end package body generics;