    -- Includes all clock generators and all sim instances (DUTs, BFMs, ...)

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;
    -- use ieee.math_complex.all;

    library std;
    use std.textio.all;
    use std.env.all;

    -- TB Packages
    --     * Module-specific TB Packages
    library lib_sim;
    use lib_sim.const_lfsr_inemul_pack_tb.all;
    use lib_sim.types_lfsr_inemul_pack_tb.all;
    use lib_sim.signals_lfsr_inemul_pack_tb.all;

    --     * Global Project-specific TB Packages
    use lib_sim.const_pack_tb.all;
    use lib_sim.types_pack_tb.all;
    use lib_sim.signals_pack_tb.all;

    --     * Generic TB Packages
    use lib_sim.print_pack_tb.all;
    use lib_sim.clk_pack_tb.all;
    use lib_sim.list_string_pack_tb.all;
    use lib_sim.print_list_pack_tb.all;

    -- SRC Packages
    --     * Module-specific SRC Packages (not used)
    -- use lib_sim.const_lfsr_inemul_pack.all;
    -- use lib_sim.types_lfsr_inemul_pack.all;
    -- use lib_sim.signals_lfsr_inemul_pack.all;

    --     * Global project-specific SRC Packages
    library lib_src;
    use lib_src.const_pack.all;
    use lib_src.types_pack.all;
    use lib_src.signals_pack.all;

    -- OSVVM Packages
    library osvvm;
    use osvvm.RandomPkg.all;


    entity harness_lfsr_inemul_tb is
    end harness_lfsr_inemul_tb;

    architecture sim of harness_lfsr_inemul_tb is
    begin

        gen_clk_freq_hz_real(clk1, real_clk1_hz);

        inst_dut_lfsr_inemul : entity lib_src.lfsr_inemul(rtl)
        port map (
            -- In
            clk => clk1,
            rst => dut1_rst,
            -- data_in  => dut1_tx1;
            -- valid_in => dut1_tx1_valid1,

            -- Out
            ready => dut1_ready,
            data_out => dut1_rx1,
            valid_out => dut1_rx1_valid1
        );


        -- DUT1 Driver: Transmit data to DUT1 on redge of clk1 if DUT1 ready
        proc_driver_dut1_tx1 : process
            variable v_dut1_tx1 : std_logic_vector(dut1_tx1'range) := (others => '0');
        begin
            if rising_edge(clk1) then
                if queue_sequence_dut1_tx1.length /= 0 then
                    if dut1_ready = '1' then
                        dut1_tx1 <= string_bits_to_slv(queue_sequence_dut1_tx1.get(0));
                        dut1_tx1_valid1 <= '1';
                    end if;
                else
                    -- dut1_tx1 <= (others => '0'); -- Uncomment for data pulldown -> monitors will have to be sensitive to dut1_tx1_valid1
                    dut1_tx1_valid1 <= '0';
                end if;
            end if;

            -- Repeat
            wait until rising_edge(clk1);
        end process;

    end architecture;