-- generics.vhd: This is an automatically generated file with generic parameters 
-- after running 'make generics' command.
package generics is

    constant INT_EMULATE_INPUTS : integer := 0;
    constant INT_QUBITS_CNT : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_1H_DELAY_NS : integer := 00;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_1H_DELAY : integer := 0;
    constant INT_ALL_DIGITS_PHOTON_1V_DELAY_NS : integer := 7;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_1V_DELAY : integer := 0;
    constant INT_ALL_DIGITS_PHOTON_2H_DELAY_NS : integer := 2046;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_2H_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_2V_DELAY_NS : integer := 2103;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_2V_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_3H_DELAY_NS : integer := 4110;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_3H_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_3V_DELAY_NS : integer := 4111;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_3V_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_4H_DELAY_NS : integer := 5773;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_4H_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_4V_DELAY_NS : integer := 5780;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_4V_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_5H_DELAY_NS : integer := -51771;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_5H_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_5V_DELAY_NS : integer := -51811;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_5V_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_6H_DELAY_NS : integer := -61771;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_6H_DELAY : integer := 3;
    constant INT_ALL_DIGITS_PHOTON_6V_DELAY_NS : integer := -61811;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_6V_DELAY : integer := 3;
    constant INT_CTRL_PULSE_HIGH_DURATION_NS : integer := 25;
    constant INT_CTRL_PULSE_DEAD_DURATION_NS : integer := 10;
    constant INT_CTRL_PULSE_EXTRA_DELAY_Q2_NS : integer := 40;
    constant INT_CTRL_PULSE_EXTRA_DELAY_Q3_NS : integer := 37;
    constant INT_CTRL_PULSE_EXTRA_DELAY_Q4_NS : integer := 2;
    constant INT_CTRL_PULSE_EXTRA_DELAY_Q5_NS : integer := 20;
    constant INT_CTRL_PULSE_EXTRA_DELAY_Q6_NS : integer := 20;
    constant INT_FEEDFWD_PROGRAMMING : integer := 01101011;

end package generics;



package body generics is 

end package body generics;