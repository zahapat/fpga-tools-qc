
    -- nff_cdcc_fedge_tb.vhd: Testbench for module nff_cdcc_fedge.vhd
    -- Engineer: Patrik Zahalka 
    -- Email: patrik.zahalka@univie.ac.at
    -- Created: 10/16/2021

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    library lib_sim;
    use lib_sim.clk_pack_tb.all;
    use lib_sim.random_pack_tb.all;

    use std.env.finish;

    library lib_src;

    entity nff_cdcc_fedge_tb is
    end nff_cdcc_fedge_tb;

    architecture sim of nff_cdcc_fedge_tb is


    begin



    end architecture;