--==========================================================================================
-- This VVC was generated with Bitvis VVC Generator
--==========================================================================================


context vvc_context is
  library vip_tx_crc_symtuppar;
  use vip_tx_crc_symtuppar.vvc_methods_pkg.all;
  use vip_tx_crc_symtuppar.td_vvc_framework_common_methods_pkg.all;
  -- use vip_tx_crc_symtuppar.tx_crc_symtuppar_bfm_pkg.t_tx_crc_symtuppar_if;
  use vip_tx_crc_symtuppar.tx_crc_symtuppar_bfm_pkg.t_tx_crc_symtuppar_bfm_config;
  use vip_tx_crc_symtuppar.tx_crc_symtuppar_bfm_pkg.C_TX_CRC_SYMTUPPAR_BFM_CONFIG_DEFAULT;
end context;
