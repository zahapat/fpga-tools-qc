
    -- memristor_ctrl_tb.vhd: Testbench for module qubit_sampler_dual_port.vhd
    -- Engineer: Patrik Zahalka 
    -- Email: patrik.zahalka@univie.ac.at
    -- Created: 10/16/2021

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    library lib_sim;
    use lib_sim.clk_pack_tb.all;
    use lib_sim.random_pack_tb.all;

    use std.env.finish;

    library lib_src;

    entity memristor_ctrl_tb is
    end memristor_ctrl_tb;

    architecture sim of memristor_ctrl_tb is



    begin



    end architecture;