    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    library lib_src;

    library lib_sim;
    use lib_sim.clk_pack_tb.all;
    use lib_sim.const_pack_tb.all;
    use lib_sim.export_pack_tb.all;
    use lib_sim.print_pack_tb.all;
    use lib_sim.random_pack_tb.all;
    use lib_sim.print_list_pack_tb.all;

    use lib_sim.list_string_pack_tb.all;

    use std.textio.all;
    use std.env.finish;
    use std.env.stop;

    entity johnson_cnt_tb is
    end johnson_cnt_tb;

    architecture sim of johnson_cnt_tb is


    begin



    end architecture;