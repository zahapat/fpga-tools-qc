    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    use std.textio.all;
    use std.env.finish;

    library lib_src;

    entity top_memristor_tb is
    end top_memristor_tb;

    architecture sim of top_memristor_tb is

        

    begin

        

    end architecture;