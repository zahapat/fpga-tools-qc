-- generics.vhd: This is an automatically generated file with generic parameters 
-- after running 'make generics' command.
package generics is

    constant INT_EMULATE_INPUTS : integer := 0;
    constant INT_QUBITS_CNT : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_1H_DELAY_NS : integer := 7565;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_1H_DELAY : integer := 2;
    constant INT_ALL_DIGITS_PHOTON_1V_DELAY_NS : integer := 7501;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_1V_DELAY : integer := 2;
    constant INT_ALL_DIGITS_PHOTON_2H_DELAY_NS : integer := -103095;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_2H_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_2V_DELAY_NS : integer := -103435;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_2V_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_3H_DELAY_NS : integer := -211735;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_3H_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_3V_DELAY_NS : integer := -212545;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_3V_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_4H_DELAY_NS : integer := -317795;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_4H_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_4V_DELAY_NS : integer := -31810;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_4V_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_5H_DELAY_NS : integer := -41771;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_5H_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_5V_DELAY_NS : integer := -41811;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_5V_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_6H_DELAY_NS : integer := -51771;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_6H_DELAY : integer := 4;
    constant INT_ALL_DIGITS_PHOTON_6V_DELAY_NS : integer := -51811;
    constant INT_WHOLE_DIGITS_CNT_PHOTON_6V_DELAY : integer := 4;
    constant INT_CTRL_PULSE_HIGH_DURATION_NS : integer := 100;
    constant INT_CTRL_PULSE_DEAD_DURATION_NS : integer := 50;
    constant INT_CTRL_PULSE_EXTRA_DELAY_NS : integer := 0;
    constant INT_DISCARD_QUBITS_TIME_NS : integer := 0;

end package generics;



package body generics is 

end package body generics;