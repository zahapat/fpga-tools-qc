    -- Constants that are accessible to all testbench modules/submodules

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

    library uvvm_util;
    context uvvm_util.uvvm_util_context;

    library uvvm_vvc_framework;
    use uvvm_vvc_framework.ti_vvc_framework_support_pkg.all;


    package const_pack_tb is

        ------------------------------------------------
        -- globally visible constants
        ------------------------------------------------
        -- USER INPUT

    end package;

    package body const_pack_tb is

    end package body;